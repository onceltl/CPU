library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.constantsIF.all;

entity TopLevel is
    Port (
		clk : in  STD_LOGIC;
		rst : in  STD_LOGIC
	);
end TopLevel;

architecture Behavioral of TopLevel is

begin


end Behavioral;

